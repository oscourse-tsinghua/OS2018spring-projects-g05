library ieee;
use ieee.std_logic_1164.all;
use work.global_const.all;

package float_const is 
end float_const;