library ieee;
use ieee.std_logic_1164.all;

package cp0_const is

    --
    -- Format of instructions, classified into R type, I type and J type
    --
    
end cp0_const;
