library ieee;
use ieee.std_logic_1164.all;
use work.global_const.all;

entity boot_ctrl is
    port (
        addr_i: in std_logic_vector(AddrWidth);
        readData_o: out std_logic_vector(DataWidth)
    );
end boot_ctrl;

architecture bhv of boot_ctrl is
    signal addr: std_logic_vector(6 downto 0);
begin
    addr <= addr_i(8 downto 2);

    with addr select readData_o <=
       "00100100000011110000000000011000" when "0011000",
       "10001101111100010000000000000000" when "0010011",
       "00000000000000000000000000000000" when "0110100",
       "00000010000011110111100000100001" when "0011001",
       "00000010000011110111100000100001" when "0010010",
       "00000000000000000000000000000000" when "0110000",
       "00100110110101100000000000000100" when "0101100",
       "00100110001100010000000000100000" when "0110001",
       "00111100000010000100011001001100" when "0001011",
       "00010010100000000000000000001100" when "0100100",
       "00100100000011110000000000101100" when "0010100",
       "00110010010100101111111111111111" when "0010111",
       "00111100000010001011111011111111" when "0000011",
       "00100100000011110000000000000000" when "0001000",
       "00000000000000000000000000000000" when "0100111",
       "10001101111101000000000000000000" when "0011101",
       "00000010000011110111100000100001" when "0100010",
       "00110101000010001111111111111000" when "0000100",
       "00000010000011110111100000100001" when "0011100",
       "00000010000011110111100000100001" when "0011111",
       "10001101111101100000000000000000" when "0100011",
       "00100110001011110000000000010000" when "0011110",
       "00010001000010010000000000000011" when "0001101",
       "10001101111100100000000000000000" when "0010110",
       "00110101000010000100010101111111" when "0001100",
       "00011110101000001111111111111000" when "0101111",
       "00000010000011110111100000100001" when "0001001",
       "00000000000000000000000000000000" when "0100101",
       "10101101000010010000000000000000" when "0000110",
       "00000000000000000000000000000000" when "0010000",
       "00100110001011110000000000001000" when "0011011",
       "00100110101101011111111111111100" when "0101110",
       "00000000000000000000000000000000" when "0111011",
       "00010000000000001111111111111111" when "0110111",
       "00000000000000000000000000000000" when "0000000",
       "00100110100101000000000000000100" when "0101101",
       "00000000000000000000000000000000" when "0110110",
       "00000000000000000000000000000000" when "0000010",
       "00010000000000000000000000000001" when "0000001",
       "00010000000000000000000000101001" when "0001111",
       "10001101111101010000000000000000" when "0100000",
       "00000000000000000000000000000000" when "0001110",
       "00100110010100101111111111111111" when "0110010",
       "00000000000000000000000000000000" when "0111000",
       "00011110010000001111111111100111" when "0110011",
       "00100110110011110000000000000000" when "0101000",
       "00111100000100001011111000000000" when "0000111",
       "00000010011000000000000000001000" when "0110101",
       "00100110001011110000000000000100" when "0100001",
       "00100100000011110000000000011100" when "0010001",
       "00000010000011110111100000100001" when "0101001",
       "00000000000000000000000000000000" when "0111010",
       "00010010101000000000000000001010" when "0100110",
       "10001101111010010000000000000000" when "0001010",
       "00010000000000001111111111111111" when "0111001",
       "10001101111010000000000000000000" when "0101010",
       "00100100000010010000000011111111" when "0000101",
       "00000010000011110111100000100001" when "0010101",
       "10001101111100110000000000000000" when "0011010",
       "10101110100010000000000000000000" when "0101011",
       "00000000000000000000000000000000" when others;
end bhv;