library ieee;
use ieee.std_logic_1164.all;
use work.global_const.all;

entity boot_ctrl is
    port (
        addr_i: in std_logic_vector(AddrWidth);
        readData_o: out std_logic_vector(DataWidth)
    );
end boot_ctrl;

architecture bhv of boot_ctrl is
    signal addr: std_logic_vector(6 downto 0);
begin
    addr <= addr_i(8 downto 2);

    with addr select readData_o <=
        "00000000000000000000000000000000" when "0000000",
        "00010000000000000000000000000001" when "0000001",
        "00000000000000000000000000000000" when "0000010",
        "00111100000010001011111011111111" when "0000011",
        "00110101000010001111111111111000" when "0000100",
        "00100100000010010000000011111111" when "0000101",
        "10101101000010010000000000000000" when "0000110",
        "00111100000100001011111000000000" when "0000111",
        "00100100000011110000000000000000" when "0001000",
        "00000010000011110111100000100001" when "0001001",
        "10001101111010010000000000000000" when "0001010",
        "10001101111011110000000000000100" when "0001011",
        "00000000000011110111110000000000" when "0001100",
        "00000001001011110100100000100101" when "0001101",
        "00111100000010000100011001001100" when "0001110",
        "00110101000010000100010101111111" when "0001111",
        "00010001000010010000000000000011" when "0010000",
        "00000000000000000000000000000000" when "0010001",
        "00010000000000000000000001000010" when "0010010",
        "00000000000000000000000000000000" when "0010011",
        "00100100000011110000000000111000" when "0010100",
        "00000010000011110111100000100001" when "0010101",
        "10001101111100010000000000000000" when "0010110",
        "10001101111011110000000000000100" when "0010111",
        "00000000000011110111110000000000" when "0011000",
        "00000010001011111000100000100101" when "0011001",
        "00100100000011110000000001011000" when "0011010",
        "00000010000011110111100000100001" when "0011011",
        "10001101111100100000000000000000" when "0011100",
        "10001101111011110000000000000100" when "0011101",
        "00000000000011110111110000000000" when "0011110",
        "00000010010011111001000000100101" when "0011111",
        "00110010010100101111111111111111" when "0100000",
        "00100100000011110000000000110000" when "0100001",
        "00000010000011110111100000100001" when "0100010",
        "10001101111100110000000000000000" when "0100011",
        "10001101111011110000000000000100" when "0100100",
        "00000000000011110111110000000000" when "0100101",
        "00000010011011111001100000100101" when "0100110",
        "00100110001011110000000000001000" when "0100111",
        "00000000000011110111100001000000" when "0101000",
        "00000010000011110111100000100001" when "0101001",
        "10001101111101000000000000000000" when "0101010",
        "10001101111011110000000000000100" when "0101011",
        "00000000000011110111110000000000" when "0101100",
        "00000010100011111010000000100101" when "0101101",
        "00100110001011110000000000010000" when "0101110",
        "00000000000011110111100001000000" when "0101111",
        "00000010000011110111100000100001" when "0110000",
        "10001101111101010000000000000000" when "0110001",
        "10001101111011110000000000000100" when "0110010",
        "00000000000011110111110000000000" when "0110011",
        "00000010101011111010100000100101" when "0110100",
        "00100110001011110000000000000100" when "0110101",
        "00000000000011110111100001000000" when "0110110",
        "00000010000011110111100000100001" when "0110111",
        "10001101111101100000000000000000" when "0111000",
        "10001101111011110000000000000100" when "0111001",
        "00000000000011110111110000000000" when "0111010",
        "00000010110011111011000000100101" when "0111011",
        "00010010100000000000000000010000" when "0111100",
        "00000000000000000000000000000000" when "0111101",
        "00010010101000000000000000001110" when "0111110",
        "00000000000000000000000000000000" when "0111111",
        "00100110110011110000000000000000" when "1000000",
        "00000000000011110111100001000000" when "1000001",
        "00000010000011110111100000100001" when "1000010",
        "10001101111010000000000000000000" when "1000011",
        "10001101111011110000000000000100" when "1000100",
        "00000000000011110111110000000000" when "1000101",
        "00000001000011110100000000100101" when "1000110",
        "10101110100010000000000000000000" when "1000111",
        "00100110110101100000000000000100" when "1001000",
        "00100110100101000000000000000100" when "1001001",
        "00100110101101011111111111111100" when "1001010",
        "00011110101000001111111111110100" when "1001011",
        "00000000000000000000000000000000" when "1001100",
        "00100110001100010000000000100000" when "1001101",
        "00100110010100101111111111111111" when "1001110",
        "00011110010000001111111111010111" when "1001111",
        "00000000000000000000000000000000" when "1010000",
        "00000010011000000000000000001000" when "1010001",
        "00000000000000000000000000000000" when "1010010",
        "00010000000000001111111111111111" when "1010011",
        "00000000000000000000000000000000" when "1010100",
        "00010000000000001111111111111111" when "1010101",
        "00000000000000000000000000000000" when "1010110",
        "00000000000000000000000000000000" when others;
end bhv;
