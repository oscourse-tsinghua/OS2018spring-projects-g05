library ieee;
use ieee.std_logic_1164.all;
use work.global_const.all;

entity boot_ctrl is
    port (
        addr_i: in std_logic_vector(AddrWidth);
        readData_o: out std_logic_vector(DataWidth)
    );
end boot_ctrl;

architecture bhv of boot_ctrl is
    signal addr: std_logic_vector(7 downto 0);
begin
    addr <= addr_i(9 downto 2);

    with addr select readData_o <=
        "00111100000000011000000000000000" when "00000000",
        "00110100001000010000000110000000" when "00000001",
        "00111100000000101011111111000000" when "00000010",
        "00110100010000100000000010001100" when "00000011",
        "00111100000000110000000001000000" when "00000100",
        "00110100011000110000000000001000" when "00000101",
        "00111100000001001011111111010000" when "00000110",
        "00110100100001000000001111111000" when "00000111",
        "00111100000001111000000000000000" when "00001000",
        "00110100111001110000001100000000" when "00001001",
        "00111100000010101000010000000000" when "00001010",
        "10101100001000110000000000000000" when "00001011",
        "10101100001000000000000000000100" when "00001100",
        "00100100000101010000000010000100" when "00001101",
        "00100100000101110111110000000001" when "00001110",
        "01000000100101110110000000000000" when "00001111",
        "00100100000110000000000000000001" when "00010000",
        "01000000100101110110000000000000" when "00010001",
        "00111100000001010000000000000100" when "00010010",
        "00100100000010000000000000000001" when "00010011",
        "00000000101010000010100000100010" when "00010100",
        "00010100101000001111111111111110" when "00010101",
        "00000000000000000000000000000000" when "00010110",
        "01000000100000000110000000000000" when "00010111",
        "00000000000000000000000000000000" when "00011000",
        "00000000000000000000000000000000" when "00011001",
        "00000000000000000000000000000000" when "00011010",
        "00000000000000000000000000000000" when "00011011",
        "00100100000001100000000000010101" when "00011100",
        "10101100111101100000000000001000" when "00011101",
        "10101100111011010000000000001100" when "00011110",
        "10101100100001100000000000000000" when "00011111",
        "00100100000101100000000000000000" when "00100000",
        "00010000000000001111111111101111" when "00100001",
        "00000000000000000000000000000000" when "00100010",
        "01000000100000000110000000000000" when "00100011",
        "00000000000000000000000000000000" when "00100100",
        "00000000000000000000000000000000" when "00100101",
        "00000000000000000000000000000000" when "00100110",
        "00000000000000000000000000000000" when "00100111",
        "10001100100011010000000000000100" when "00101000",
        "00100100000000110000000000000010" when "00101001",
        "00010001101000110000000000000110" when "00101010",
        "00000000000000000000000000000000" when "00101011",
        "00100100000000110000000000000011" when "00101100",
        "00010001101000110000000000000011" when "00101101",
        "00000000000000000000000000000000" when "00101110",
        "00010000000000001111111111100001" when "00101111",
        "00000000000000000000000000000000" when "00110000",
        "00100110110101100000000000000001" when "00110001",
        "10001100100011010000000000000000" when "00110010",
        "00100100000000110000000000000001" when "00110011",
        "00010010110000110000000000011010" when "00110100",
        "00000000000000000000000000000000" when "00110101",
        "00100100000000110000000000000010" when "00110110",
        "00010010110000110000000000011111" when "00110111",
        "00000000000000000000000000000000" when "00111000",
        "00100100000000110000000000000011" when "00111001",
        "00010010110000110000000000100011" when "00111010",
        "00000000000000000000000000000000" when "00111011",
        "00100100000000110000000000000100" when "00111100",
        "00000010110000110001100000100011" when "00111101",
        "00000000111000111100100000100000" when "00111110",
        "00100100000110100000000000000011" when "00111111",
        "00000011010110011101100000100100" when "01000000",
        "00000011001110111110000000100010" when "01000001",
        "10001111100110100000000000000000" when "01000010",
        "00100100000110010000000011111111" when "01000011",
        "00000000000110111101100011000000" when "01000100",
        "00000011011110011100100000000100" when "01000101",
        "00000011001110101100100000100100" when "01000110",
        "00000011010110011101000000100110" when "01000111",
        "00000011011011011101100000000100" when "01001000",
        "00000011010110111101000000100000" when "01001001",
        "10101111100110100000000000000000" when "01001010",
        "00010010110101010000000000011000" when "01001011",
        "00000000000000000000000000000000" when "01001100",
        "00010000000000001111111111000011" when "01001101",
        "00000000000000000000000000000000" when "01001110",
        "00100100000000110000000000000100" when "01001111",
        "00010001101000110000000001000101" when "01010000",
        "00000000000000000000000000000000" when "01010001",
        "00100100000000110000000000000001" when "01010010",
        "00010001101000111111111110111101" when "01010011",
        "00000000000000000000000000000000" when "01010100",
        "00010000000000001111111111000110" when "01010101",
        "00000000000000000000000000000000" when "01010110",
        "00100101101101000000000000000001" when "01010111",
        "00010010100110000000000000110110" when "01011000",
        "00000000000000000000000000000000" when "01011001",
        "00010001101110001111111110110110" when "01011010",
        "00000000000000000000000000000000" when "01011011",
        "00010000000000001111111110111111" when "01011100",
        "00000000000000000000000000000000" when "01011101",
        "00100100000000110000000011111111" when "01011110",
        "00000000011110000001100000100011" when "01011111",
        "00010000011011011111111110110000" when "01100000",
        "00000000000000000000000000000000" when "01100001",
        "00010000000000001111111110111001" when "01100010",
        "00000000000000000000000000000000" when "01100011",
        "00100100000010110000000010000000" when "01100100",
        "00100100000011000000000000000000" when "01100101",
        "00100100000011010000000000000000" when "01100110",
        "00000000111011001100100000100000" when "01100111",
        "00100100000110100000000000000011" when "01101000",
        "00000011010110011101100000100100" when "01101001",
        "00000011001110111110000000100010" when "01101010",
        "10001111100110100000000000000000" when "01101011",
        "00100100000110010000000011111111" when "01101100",
        "00000000000110111101100011000000" when "01101101",
        "00000011011110011100100000000100" when "01101110",
        "00000011010110011101000000100100" when "01101111",
        "00000011011110100111000000000110" when "01110000",
        "00100101100011000000000000000001" when "01110001",
        "00000001101011100110100000100000" when "01110010",
        "00010101100010111111111111110011" when "01110011",
        "00000000000000000000000000000000" when "01110100",
        "00110001101011010000000011111111" when "01110101",
        "00000000111011001100100000100000" when "01110110",
        "00100100000110100000000000000011" when "01110111",
        "00000011010110011101100000100100" when "01111000",
        "00000011001110111110000000100010" when "01111001",
        "10001111100110100000000000000000" when "01111010",
        "00100100000110010000000011111111" when "01111011",
        "00000000000110111101100011000000" when "01111100",
        "00000011011110011100100000000100" when "01111101",
        "00000011010110011101000000100100" when "01111110",
        "00000011011110100111000000000110" when "01111111",
        "00100101100011000000000000000001" when "10000000",
        "00010001101011100000000000000011" when "10000001",
        "00000000000000000000000000000000" when "10000010",
        "00010000000000001111111110011000" when "10000011",
        "00000000000000000000000000000000" when "10000100",
        "00100100000010110000000000000000" when "10000101",
        "00100100000011000000000000100000" when "10000110",
        "00000000111000000110100000100101" when "10000111",
        "00100101101011010000000000000100" when "10001000",
        "00100101010010100000000000000100" when "10001001",
        "10001101101011101111111111111100" when "10001010",
        "10101101010011101111111111111100" when "10001011",
        "00100101011010110000000000000001" when "10001100",
        "00010101011011001111111111111010" when "10001101",
        "00000000000000000000000000000000" when "10001110",
        "00100100000001100000000000000110" when "10001111",
        "10101100100001100000000000000000" when "10010000",
        "00100100000101100000000000000000" when "10010001",
        "00100111000110000000000000000001" when "10010010",
        "00110011000110000000000011111111" when "10010011",
        "00010000000000001111111101111100" when "10010100",
        "00000000000000000000000000000000" when "10010101",
        "00100100000001100000000000000110" when "10010110",
        "10101100100001100000000000000000" when "10010111",
        "01000000100000000110000000000000" when "10011000",
        "00111100000010001000011111111111" when "10011001",
        "00110101000010001111111111111000" when "10011010",
        "00100100000010010000000011111111" when "10011011",
        "10101101000010010000000000000000" when "10011100",
        "00111100000100001000010000000000" when "10011101",
        "00100100000011110000000000000000" when "10011110",
        "00000010000011110111100000100001" when "10011111",
        "10001101111010010000000000000000" when "10100000",
        "00111100000010000100011001001100" when "10100001",
        "00110101000010000100010101111111" when "10100010",
        "00010001000010010000000000000011" when "10100011",
        "00000000000000000000000000000000" when "10100100",
        "00010000000000000000000000100111" when "10100101",
        "00000000000000000000000000000000" when "10100110",
        "00100100000011110000000000011100" when "10100111",
        "00000010000011110111100000100001" when "10101000",
        "10001101111100010000000000000000" when "10101001",
        "00100100000011110000000000101100" when "10101010",
        "00000010000011110111100000100001" when "10101011",
        "10001101111100100000000000000000" when "10101100",
        "00110010010100101111111111111111" when "10101101",
        "00100100000011110000000000011000" when "10101110",
        "00000010000011110111100000100001" when "10101111",
        "10001101111100110000000000000000" when "10110000",
        "00100110001011110000000000001000" when "10110001",
        "00000010000011110111100000100001" when "10110010",
        "10001101111101000000000000000000" when "10110011",
        "00100110001011110000000000010000" when "10110100",
        "00000010000011110111100000100001" when "10110101",
        "10001101111101010000000000000000" when "10110110",
        "00100110001011110000000000000100" when "10110111",
        "00000010000011110111100000100001" when "10111000",
        "10001101111101100000000000000000" when "10111001",
        "00010010100000000000000000001100" when "10111010",
        "00000000000000000000000000000000" when "10111011",
        "00010010101000000000000000001010" when "10111100",
        "00000000000000000000000000000000" when "10111101",
        "00100110110011110000000000000000" when "10111110",
        "00000010000011110111100000100001" when "10111111",
        "10001101111010000000000000000000" when "11000000",
        "10101110100010000000000000000000" when "11000001",
        "00100110110101100000000000000100" when "11000010",
        "00100110100101000000000000000100" when "11000011",
        "00100110101101011111111111111100" when "11000100",
        "00011110101000001111111111111000" when "11000101",
        "00000000000000000000000000000000" when "11000110",
        "00100110001100010000000000100000" when "11000111",
        "00100110010100101111111111111111" when "11001000",
        "00011110010000001111111111100111" when "11001001",
        "00000000000000000000000000000000" when "11001010",
        "00000010011000000000000000001000" when "11001011",
        "00000000000000000000000000000000" when "11001100",
        "00010000000000001111111111111111" when "11001101",
        "00000000000000000000000000000000" when "11001110",
        "00000000000000000000000000000000" when "11001111",
        "00000000000000000000000000000000" when others;
end bhv;
